module sdio_device_phy_sd_ls (
  input               clk,
  input               rst,

  //PHY Layer
  output              ddr_en,
  input               sdio_clk,
  input               sdio_cs_n,
  input [3:0]         sdio_data


);
//Local Parameters

//Local Registers/Wires
//Submodules


//Asynchronous Logic
//Synchronous Logic


endmodule


